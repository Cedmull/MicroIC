library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

package sprite_book is
    type sprite is array (natural range 0 to 2499) of std_logic_vector(11 downto 0);
    constant red_square : sprite := ( "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011", "111001000011");
    constant blue_square : sprite := ( "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101", "001110011101");
end sprite_book;