package sprite_book is
    type sprite is array (natural range 0 to 2499) of std_logic_vector(11 downto 0);
    constant red_square : sprite := ( "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110", "111011101110");
    constant blue_square : sprite := ( "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011", "001100110011");
end sprite_book;
